// Register group