// Register group
module regs(
    input logic clk,
    input logic [4:0] 
)