    //============================
    //        FSM for AXI
    //============================